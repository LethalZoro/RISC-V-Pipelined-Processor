module tb;
wire  ;
reg  ;

top uut(
    .(),
    .(),
    .()
);

initial begin

    #100;
end

endmodule